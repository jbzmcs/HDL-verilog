module notGate_df(input a, output b);
    assign b = ~a;
endmodule