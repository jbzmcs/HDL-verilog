module notGate_st(input a, output b);
    not not1(b,a);
endmodule