module and(a,b);
    input a,b;
    output y;

    //and (a,b);
    assign y = a + b;

endmodule