module xorGate_df(input a,b, output c);
    assign c = a ^ b; // xor operator
endmodule