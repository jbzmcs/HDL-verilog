//Structural
module orGateLab1_st(input wire a,b, output wire c);
    or or1(c,a,b);
    
endmodule